module hardware

